// FPGA Top Level

`default_nettype none

module top (
 // I/O ports
  input  logic hz100, reset,
  input  logic [20:0] pb,
  output logic [7:0] left, right,
         ss7, ss6, ss5, ss4, ss3, ss2, ss1, ss0,
  output logic red, green, blue,

  // UART ports
  output logic [7:0] txdata,
  input  logic [7:0] rxdata,
  output logic txclk, rxclk,
  input  logic txready, rxready

);
// assign right [0] = 1'b1;
logic [31:0] display;
top1 top (.clk(pb[18]), .nrst(!pb[19]), .display(display));
ssdec s7 (.in(display[15:12]), .enable(1'b1), .out(ss7[6:0]));
ssdec s6 (.in(display[11:8]), .enable(1'b1), .out(ss6[6:0]));
ssdec s5 (.in(display[7:4]), .enable(1'b1), .out(ss5[6:0]));
ssdec s4 (.in(display[3:0]), .enable(1'b1), .out(ss4[6:0]));



endmodule
